*DIODES_INC_SPICE_MODEL
*ORIGIN=DZSL_DPG_GM
*SIMULATOR=PSPICE
*DATE=08FEB2011
*VERSION=2
*
.MODEL MMBT5551 NPN IS=6.5E-15 NF=1 BF=110 VAF=288 ISE=1.0E-14
+ NE=1.5 NR=1 BR=4.5 VAR=70 ISC=3E-12 NC=1.35 RC=0.5 RB =0.26 RE =0.23
+ CJC=6.1E-12 MJC=0.31 VJC=0.4 CJE=57E-12 MJE=0.35 VJE=0.8 TF=0.2E-9
+ TR=1.5E-6 XTB=1.4 QUASIMOD=1 RCO=170 VO=35 GAMMA=2.2E-7
*
*$
