*---------- 5N10 MOSFET SPICE Model (Chatgpt generated) ----------
.SUBCKT 5N10 D G S
*     TERMINALS:  D  G  S
M1 D G S S NMOS L=1E-006 W=50E-006
RD D Dint 0.12
RS S Sint 0.01
RG G Gint 10
CGS G S 1.2E-10
CGD G D 3.5E-11
.MODEL NMOS NMOS LEVEL=3 VTO=2 KP=120 U0=600 VMAX=5E5
+ TOX=8E-008 NSUB=1E16 KAPPA=10
.MODEL Dint D IS=1E-12 BV=100 CJO=3E-12 VJ=0.7 M=0.5
.MODEL Sint D IS=1E-12
.ENDS
