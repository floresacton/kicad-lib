*---------- BSS123(Z) Spice Model ----------
.SUBCKT BSS123Z 10 20 30 
*     TERMINALS:  D  G  S
M1 1 2 3 3 NMOS L = 1E-006 W = 1E-006 
RD 10 1 2.298 
RS 30 3 0.001 
RG 20 2 17 
CGS 2 3 5.7E-011 
EGD 12 0 2 1 1 
VFB 14 0 0 
FFB 2 1 VFB 1 
CGD 13 14 1E-011 
R1 13 0 1 
D1 12 13 DLIM 
DDG 15 14 DCGD 
R2 12 15 1 
D2 15 0 DLIM 
DSD 3 10 DSUB 
.MODEL NMOS NMOS LEVEL = 3 VMAX = 5.378E+005 ETA = 0.001 VTO = 1.75 
+ TOX = 6E-008 NSUB = 1E+016 KP = 1.58 U0 = 400 KAPPA = 10 
.MODEL DCGD D CJO = 1.2E-011 VJ = 0.8 M = 0.6 
.MODEL DSUB D IS = 1.847E-009 N = 1.638 RS = 0.1103 BV = 115 CJO = 1E-011 VJ = 0.7586 M = 0.6096 
.MODEL DLIM D IS = 0.0001 
.ENDS
*Diodes BSS123Z Spice Model v1.0M Last Revised 2016/10/6
